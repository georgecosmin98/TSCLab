/***********************************************************************
 * A SystemVerilog testbench for an instruction register; This file
 * contains the interface to connect the testbench to the design
 *
 * SystemVerilog Training Workshop.
 * Copyright 2006, 2013 by Sutherland HDL, Inc.
 * Tualatin, Oregon, USA.  All rights reserved.
 * www.sutherland-hdl.com
 **********************************************************************/
interface tb_ifc (input logic clk);
  timeunit 1ns/1ns;

  // user-defined types are defined in instr_register_pkg.sv
  import instr_register_pkg::*;

  // ADD CODE TO DECLARE THE INTERFACE SIGNALS
  logic          load_en; 
  logic          reset_n;
  opcode_t       opcode;
  operand_t      operand_a, operand_b;
  address_t      write_pointer, read_pointer;
  instruction_t  instruction_word;

  // ADD CODE TO DEFINE A CLOCKING BLOCK WITH INPUT AND OUTPUT SKEWS
  clocking cb @(posedge clk); //declare cb
    output load_en;
    output reset_n;
    output opcode;
    output operand_a;
    output operand_b;
    output write_pointer;
    output read_pointer;
    input instruction_word;
  endclocking

  //modport TEST (clocking cb);

 // modport DUT (input load_en,
  //             input reset_n,
 //              input opcode,
  //             input operand_a,
 //              input operand_b,
 //              input write_pointer,
 //              input read_pointer,
 //              input instruction_word);

endinterface: tb_ifc

